library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package de2_115_seven_segment is
	type SEG_ARR is array(0 TO 7) of std_logic_vector(6 downto 0);
end package;

package body de2_115_seven_segment is
end de2_115_seven_segment;